--
-- VHDL Architecture ece411.Test1.untitled
--
-- Created:
--          by - adalton2.ews (gelib-057-31.ews.illinois.edu)
--          at - 21:12:27 02/13/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY Test1 IS
-- Declarations

END Test1 ;

--
ARCHITECTURE untitled OF Test1 IS
BEGIN
END ARCHITECTURE untitled;

